//Legal Notice: (C)2007 Altera Corporation. All rights reserved.  Your
//use of Altera Corporation's design tools, logic functions and other
//software and tools, and its AMPP partner logic functions, and any
//output files any of the foregoing (including device programming or
//simulation files), and any associated documentation or information are
//expressly subject to the terms and conditions of the Altera Program
//License Subscription Agreement or other applicable license agreement,
//including, without limitation, that your use is for the sole purpose
//of programming logic devices manufactured by Altera and sold by Altera
//or its authorized distributors.  Please refer to the applicable
//agreement for further details.

// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module Double_ADS805_0 (
                         // inputs:
                          ad_clk,
                          address,
                          clk,
                          i_input,
                          read,
                          rst_n,
                          u_input,
                          write,
                          writedata,

                         // outputs:
                          irq,
                          readdata
                       )
;

  output           irq;
  output  [ 31: 0] readdata;
  input            ad_clk;
  input   [  1: 0] address;
  input            clk;
  input   [ 11: 0] i_input;
  input            read;
  input            rst_n;
  input   [ 11: 0] u_input;
  input            write;
  input   [ 31: 0] writedata;

  wire             irq;
  wire    [ 31: 0] readdata;
  Double_ADS805 the_Double_ADS805
    (
      .ad_clk    (ad_clk),
      .address   (address),
      .clk       (clk),
      .i_input   (i_input),
      .irq       (irq),
      .read      (read),
      .readdata  (readdata),
      .rst_n     (rst_n),
      .u_input   (u_input),
      .write     (write),
      .writedata (writedata)
    );


endmodule

